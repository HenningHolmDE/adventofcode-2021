entity day_01 is
end entity;

architecture simulation of day_01 is

begin

    process
    begin
        report "Hello, world!";
        wait;
    end process;

end architecture;